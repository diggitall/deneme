module git_test_module(
    input   i_inp_1,
    input   i_inp_2,
    output  o_outp_1
  );
  
  // Test module
  
endmodule